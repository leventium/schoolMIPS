`define GPIO_SIZE 16
